library ieee;
use ieee.std_logic_1164.all;

entity SR is
	port(A: in std_logic_vector(15 downto 0);
	output: out std_logic_vector(15 downto 0));
end SR ;

architecture SR of SR is
begin
	output <= '0' & A(15 downto 1);
end SR;